`ifndef CFS_ALGN_TEST_PKG_SV
    `define CFS_ALGN_TEST_PKG_SV
package cfs_algn_test_pkg;
  
    `include "cfs_algn_test_base.sv"
    `include "cfs_algn_test_reg_access.sv"

endpackage : cfs_algn_test_pkg

`endif // CFS_ALGN_TEST_PKG_SV